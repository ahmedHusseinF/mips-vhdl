library ieee ;
  use ieee.std_logic_1164.all ;
  use ieee.numeric_std.all ;

entity cpu is
  port (
    clock: in std_logic
  );
end cpu; 

architecture cpu_wiring of cpu is

begin

  -- to implement

end architecture;