library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity cpu_test is
  generic (n: integer := 16);
end cpu_test;


architecture cpu_test_arch of cpu_test is

begin


end cpu_test_arch; -- ImpTestBench